"Unknown testcase circuit10