"Unknown testcase clock