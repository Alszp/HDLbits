"Unknown testcase ece241_2014_q4