"Unknown testcase circuit2