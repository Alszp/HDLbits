"Unknown testcase circuit5