module top_module(
    input [31:0] a,
    input [31:0] b,
    output [31:0] sum
);
    wire carryout;
    add16 numbah1(a[15:0],b[15:0],,sum[15:0],carryout);
    add16 numbah2(a[31:16],b[31:16],carryout,sum[31:16]);
endmodule
