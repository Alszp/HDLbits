"Unknown testcase tb2