"Unknown testcase review2015_fsmonehot