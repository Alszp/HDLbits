"Unknown testcase review2015_fsm