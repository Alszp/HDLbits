"Unknown testcase 2014_q4a