"Unknown testcase ece241_2013_q8