"Unknown testcase 2014_q3fsm