"Unknown testcase m2014_q4c