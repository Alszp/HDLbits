"Unknown testcase circuit1