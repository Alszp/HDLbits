"Unknown testcase circuit6