"Unknown testcase circuit8