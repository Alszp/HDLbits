"Unknown testcase m2014_q3