"Unknown testcase review2015_shiftcount