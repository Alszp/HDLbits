"Unknown testcase and