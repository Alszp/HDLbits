"Unknown testcase review2015_count1k