"Unknown testcase tff