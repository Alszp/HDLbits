"Unknown testcase 2012_q1g