"Unknown testcase circuit7