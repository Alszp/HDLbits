"Unknown testcase circuit9