"Unknown testcase circuit3