"Unknown testcase review2015_fsmshift