"Unknown testcase tb1