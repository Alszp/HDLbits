"Unknown testcase review2015_fancytimer