"Unknown testcase review2015_fsmseq