"Unknown testcase circuit4