"Unknown testcase m2014_q4h